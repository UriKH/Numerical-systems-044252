// Smart traffic system testbench
module traffic_system_smart(
    input logic clk,
    input logic reset,
    input logic start,
    input logic person_present,
    input logic car_present,
    output logic [1:0] L_out
);

// Enter X and Y here
	localparam X = 1;
	localparam Y = 2;

// Put your code here
// ------------------


// End of your code
endmodule
