// 32X32 Multiplier test template
module traffic_system(
    input logic clk,
    input logic reset,
    input logic start,
    output logic [1:0] L_out
);

// Enter X and Y here
	localparam X = 1;
	localparam Y = 2;

// Put your code here
// ------------------


// end of your code
endmodule
