// Smart timer module

module timer_smart(
    input logic clk,
    input logic reset,
    input logic t_start,
    input logic[4:0] t_length,
    input logic t_freeze,

    output logic t_flicker,
    output logic t_done
);

// Put your code here
// ------------------

//end of your code
endmodule